`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/12/2022 10:30:32 PM
// Design Name: 
// Module Name: Instruction_Memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Instruction_Memory(read_addr, instruction, reset);
input reset;
input [7:0] read_addr;
output [31:0] instruction;
reg [31:0] Imemory [63:0];
integer k;
// I-MEM in this case is addressed by word, not by byte
wire [5:0] shifted_read_addr;
assign shifted_read_addr=read_addr[7:2];
assign instruction = Imemory[shifted_read_addr];
always @(posedge reset)
begin
    for (k=30; k<64; k=k+1) begin// here Ou changes k=0 to k=16
    Imemory[k] = 32'b0;
    end
    Imemory[0] = 32'b10001101000010000000000000000000; //lw $t0,0($0)
    Imemory[1] = 32'b10001101000010010000000000000001; //lw $t1,1($0)
    Imemory[2] = 32'b10001101000010100000000000000010; //lw $t2,2($0)
    Imemory[3] = 32'b10001101000010110000000000000011; //lw $t3,3($0)
    Imemory[4] = 32'b10001101000011000000000000000100; //lw $t4,4($0)
    
    Imemory[5] = 32'b10001101000010000000000000000000; //lw $t0,0($0)
    Imemory[6] = 32'b10001101000010010000000000000001; //lw $t1,1($0)
    Imemory[7] = 32'b10001101000010100000000000000010; //lw $t2,2($0)
    Imemory[8] = 32'b10001101000010110000000000000011; //lw $t3,3($0)
    Imemory[9] = 32'b10001101000011000000000000000100; //lw $t4,4($0)
    Imemory[10] = 32'b10101101000010000000000000011111; //sw $t0,31($0)
    Imemory[11] = 32'b10101101000010010000000000100000; //sw $t1,32($0)
    Imemory[12] = 32'b10101101000010100000000000100001; //sw $t2,33($0)
    Imemory[13] = 32'b10101101000010110000000000100010; //sw $t3,34($0)
    Imemory[14] = 32'b10101101000011000000000000100011; //sw $t4,35($0)
    
    Imemory[15] = 32'b10001101000010000000000000000000; //lw $t0,0($0)
    Imemory[16] = 32'b10001101000010010000000000000001; //lw $t1,1($0)
    Imemory[17] = 32'b10001101000010100000000000000010; //lw $t2,2($0)
    Imemory[18] = 32'b10001101000010110000000000000011; //lw $t3,3($0)
    Imemory[19] = 32'b10001101000011000000000000000100; //lw $t4,4($0)
    Imemory[20] = 32'b00000001000011001000000000100000; //add $s0, $t0,$t4
    Imemory[21] = 32'b00000010000011001000100000100010; //sub $s1,$s0,$t4
    Imemory[22] = 32'b00000001010100011001000000100000; //add $s2,$t2,$s1
    Imemory[23] = 32'b00010010000100110000000000001010; //SLL $s3,$s2,4
    Imemory[24] = 32'b10101101000100000000000000100000; //SW $s0, 32($0)
    Imemory[25] = 32'b10101101100111000111111111111111; //SW $s1, -1($s3)
    
    Imemory[26] = 32'b00100000000001010110100000010000; //addi $t5, $0,5
    Imemory[27] = 32'b00100001101111010111000000010000; //addi $t6,$t5,-3
    Imemory[28] = 32'b10001101000010000000000000000000; //lw $t0,0($0)
    Imemory[29] = 32'b10001101000010010000000000000001; //lw $t1,1($0)
    Imemory[30] = 32'b10001101000010100000000000000010; //lw $t2,2($0)
    Imemory[31] = 32'b10001101000010110000000000000011; //lw $t3,3($0)
    Imemory[32] = 32'b10001101000011000000000000000100; //lw $t4,4($0)
    Imemory[33] = 32'b00000001000011001000000000100000; //add $s0,$t0,$t4
    Imemory[34] = 32'b00000010000011001000100000100010; //sub $s1,$s0,$t4
    Imemory[35] = 32'b00000001010100011001000000100000; //add $s2,$s1,$t2
    end
endmodule
