`timescale 1ns / 1ps

module MEM(    
    input clk,
    input MWE,
    input [31:0] MRA,
    input [31:0] MWD,
    output [31:0] MRD
    );
    
    reg [31:0] Memory [550:0]; // 32-bit memory
    
    initial begin
        // Memory Values
        Memory[0] <= 17; // h'00000011
        Memory[1] <= 31; // h'00000000
        Memory[2] <= -5; // h'00000000
        Memory[3] <= -2; // h'00000000
        Memory[4] <= 250; // h'00000000
        
        // PART A
//        Memory[500] <= 32'b10001100000010000000000000000000; // LW $t0 0($0) (h'8C080000)
//        Memory[501] <= 32'b10001100000010010000000000000001; // LW $t1 1($0) (h'8C090001)
//        Memory[502] <= 32'b10001100000010100000000000000010; // LW $t2 2($0) (h'8C0A0002)
//        Memory[503] <= 32'b10001100000010110000000000000011; // LW $t3 3($0) (h'8C0B0003)
//        Memory[504] <= 32'b10001100000011000000000000000100; // LW $t4 4($0) (h'8C0C0004)

//         PART B
//        Memory[500] <= 32'b10001100000010000000000000000000; // LW $t0 0($0) (h'8C080000)
//        Memory[501] <= 32'b10001100000010010000000000000001; // LW $t1 1($0) (h'8C090001)
//        Memory[502] <= 32'b10001100000010100000000000000010; // LW $t2 2($0) (h'8C0A0002)
//        Memory[503] <= 32'b10001100000010110000000000000011; // LW $t3 3($0) (h'8C0B0003)
//        Memory[504] <= 32'b10001100000011000000000000000100; // LW $t4 4($0) (h'8C0C0004)
//        Memory[505] <= 32'b10101100000010000000000000011111; // SW $t0 31($0)
//        Memory[506] <= 32'b10101100000010010000000000100000; // SW $t1 32($0)
//        Memory[507] <= 32'b10101100000010100000000000100001; // SW $t2 33($0)
//        Memory[508] <= 32'b10101100000010110000000000100010; // SW $t3 34($0)
//        Memory[509] <= 32'b10101100000011000000000000100011; // SW $t4 35($0)
       
        // PART C
//        Memory[500] <= 32'b10001100000010000000000000000000; // LW $t0 0($0) (h'8C080000)
//        Memory[501] <= 32'b10001100000010010000000000000001; // LW $t1 1($0) (h'8C090001)
//        Memory[502] <= 32'b10001100000010100000000000000010; // LW $t2 2($0) (h'8C0A0002)
//        Memory[503] <= 32'b10001100000010110000000000000011; // LW $t3 3($0) (h'8C0B0003)
//        Memory[504] <= 32'b10001100000011000000000000000100; // LW $t4 4($0) (h'8C0C0004)
//        Memory[505] <= 32'b00000001000011001000000000100000; // ADD $s0, $t0, $t4
//        Memory[506] <= 32'b00000010000011001000100000100010; // SUB $s1, $s0, $t4
//        Memory[507] <= 32'b00000001010100011001000000100000; // ADD $s2, $t2, $s1
//        Memory[508] <= 32'b00000000000100101001100100000000; // SLL $s3, $s2, 4
//        Memory[509] <= 32'b10101100000100000000000000100000; // SW $s0, 32($0)
//        Memory[510] <= 32'b10101110011100011111111111111111; // SW $s1, -1($s0)
        
        // PART D
//        Memory[500] <= 32'b00100000000011010000000000000101; // ADDI $t5, $0, 5
//        Memory[501] <= 32'b00100001101011101111111111111101; // ADDI $t6, $t5, -3      
//        Memory[502] <= 32'b10001100000010000000000000000000; // LW $t0 0($0) (h'8C080000)
//        Memory[503] <= 32'b10001100000010010000000000000001; // LW $t1 1($0) (h'8C090001)
//        Memory[504] <= 32'b10001100000010100000000000000010; // LW $t2 2($0) (h'8C0A0002)
//        Memory[505] <= 32'b10001100000010110000000000000011; // LW $t3 3($0) (h'8C0B0003)
//        Memory[506] <= 32'b10001100000011000000000000000100; // LW $t4 4($0) (h'8C0C0004)      
//        Memory[507] <= 32'b00000001000011001000000000100000; // ADD $s0, $t0, $t4
//        Memory[508] <= 32'b00000010000011001000100000100010; // SUB $s1, $s0, $t4
//        Memory[509] <= 32'b00000001010100011001000000100000; // ADD $s2, $t2, $s1             
//        Memory[510] <= 32'b00000001101100101001100000000100; // SLLV $s3, $s2, $t5
//        Memory[511] <= 32'b00000001110100101010000000000111; // SRAV $s4, $s2, $t6
//        Memory[512] <= 32'b10101100000100000000000000100000; // SW $s0, 32($0)
//        Memory[513] <= 32'b10101110011100010000000000000000; // SW $s1, 0($s3)
//        Memory[514] <= 32'b10101110100100010000000000000000; // SW $s1, 0($s4)
        
        // PART E
        Memory[500] <= 32'b00100000000100000000000000000000; // ADDI $s0, $0, 0
        Memory[501] <= 32'b00100000000100010000000000000101; // ADDI $s1, $0, 5
        Memory[502] <= 32'b00100000000100100000000000000001; // ADDI $s2, $0, 1
        Memory[503] <= 32'b00000000000000000101100000100000; // ADD $t3, $0, $0
        Memory[504] <= 32'b00010010000100010000000000000110; // loop: BEQ $s0, $s1, done
        Memory[505] <= 32'b10001110000010000000000000000000; // LW $t0, 0($s0)
        Memory[506] <= 32'b00000010001010000100000000000100; // SLLV $t0, $t0, $s1
        Memory[507] <= 32'b10101110000010000000000000011111; // SW $t0, 31($s0)
        Memory[508] <= 32'b00000010010100001000000000100000; // ADD $s0, $s2, $s
        Memory[509] <= 32'b00000001011010000101100000100000; // ADD $t3, $t3, $t
        Memory[510] <= 32'b00001000000000001111111111111001; // J loop
        Memory[511] <= 32'b00000000000000000000000000100000; // done: NOP (add $0, $0, $0)
        Memory[512] <= 32'b00000000000000000000000000100000; // NOP (add $0, $0, $0)
    end
    
    assign MRD = Memory[MRA];
    
    always@(posedge clk) begin
        if (MWE) begin
            Memory[MRA] <= MWD; // Write data DMWD onto address DMA 
        end
    end
endmodule
